module mux7sig(
  input  logic clk,
  input  logic reset,
  input  logic[15:0] switch,
  input  logic[11:0] led,
  output logic[7:0] an,
  output logic[6:0] a2g
);

endmodule